
// ???? Verilog
// ????? ???'?????? ?????
// ????????: ???? 3 - Testbench ??? spi_master

// ???????????? ??????? ????: 1?? = ???? ?????????, 1?? = ????????
`timescale 1ns / 1ps 

// ??? ?????? ????????? ?? ??? ??????, ??? "????" ??? ? ????
module spi_tb;

    /* --- ????????? ????????? --- */
    localparam CLK_PERIOD = 10; // ?????? CLK = 10?? (100???)

    /* --- ??????? ??? ??????????? ?? ?????? ?????? (DUT) --- */
    // 'reg' - ?? ???????, ????? ????? ??? testbench (????? ??????)
    reg        tb_clk;       
    reg        tb_rst_n;     
    reg        tb_start_tx;  
    reg  [7:0] tb_tx_data;   
    reg        tb_miso;      // ?? ???????? Slave, ???? ?? 'reg'
    
    // 'wire' - ?? ???????, ??? ??????? ??? ?????? (?????? ??????)
    wire       tb_tx_done;   
    wire [7:0] tb_rx_data;   
    wire       tb_sck;       
    wire       tb_mosi;      
    wire       tb_ss;        

    /* --- 1. "?????????" ?????? ?????? (DUT - Device Under Test) --- */
    // ??? ?? "??????????" ??? spi_master ? ??? ????????
    // ? ??????????? ???? 'reg' ?? 'wire' ?? ???? ??????
    spi_master DUT (
        .i_clk(tb_clk),
        .i_rst_n(tb_rst_n),
        .i_start_tx(tb_start_tx),
        .i_tx_data(tb_tx_data),
        .o_tx_done(tb_tx_done),
        .o_rx_data(tb_rx_data),
        .o_sck(tb_sck),
        .o_mosi(tb_mosi),
        .i_miso(tb_miso),
        .o_ss(tb_ss)
    );

    /* --- 2. ????????? CLK --- */
    // ??? ???? 'initial' ??????????? ???? ??? ?? ???????
    // ? ??????? ???????? ?????? ??????????? 
    initial begin
        tb_clk = 0;
        forever #(CLK_PERIOD / 2) tb_clk = ~tb_clk;
    end

    /* --- 3. ???????? Slave-???????? (????? MISO) --- */
    // ??? ???? ?????? ????????? Slave-????????.
    // ??? ??????, ?? Master (??? ??????) ????? ?????????? (tb_ss ???? 0)
    // ? ?? ????? ???? SCK ?????????? ????? ?????? ???? (??? - 8'hAA)
    reg [7:0] slave_shift_reg;
    always @(negedge tb_ss or posedge tb_sck) begin
        if (!tb_ss) begin 
            // ?? ?????? SS ???????????, ???????????? ???? ??? ?????????
            slave_shift_reg <= 8'hAA; // ?????????? ???? 10101010
        end
        
        // (CPHA=0): Slave ????????? ???? ??? ?? negedge SCK
        if (!tb_ss && tb_sck == 0) begin
            tb_miso <= slave_shift_reg[7];
            slave_shift_reg <= {slave_shift_reg[6:0], 1'b0};
        end
    end

    /* --- 4. ???????? ????????? (Test Case) --- */
    // ??? ???? 'initial' ??????, ?? ??? ???????????
    // ----- ????? ??? (?????????) -----
// ----- ????? ??? (?????????) -----
initial begin
    $display("Simulation Started..."); // <-- ???????
    // 1) ???????? ???????
    tb_rst_n = 0; 
    tb_start_tx = 0;
    tb_tx_data = 8'd0;
    #(CLK_PERIOD * 3); 
    tb_rst_n = 1; 
    #(CLK_PERIOD);

    // 2) ???????? ??????? 1: ????????? 0x55
    $display("Test 1: Sending 0x55..."); // <-- ???????
    tb_tx_data = 8'h55; 
    tb_start_tx = 1; 
    #(CLK_PERIOD);
    tb_start_tx = 0; 

    wait (tb_tx_done == 1);
    $display("Test 1 Complete. Received: %h", tb_rx_data); // <-- ???????
    #(CLK_PERIOD * 5); 

    // 3) ???????? ??????? 2: ????????? 0xF0
    $display("Test 2: Sending 0xF0..."); // <-- ???????
    tb_tx_data = 8'hF0; 
    tb_start_tx = 1;
    #(CLK_PERIOD);
    tb_start_tx = 0;

    wait (tb_tx_done == 1);
    $display("Test 2 Complete. Received: %h", tb_rx_data); // <-- ???????
    #(CLK_PERIOD * 5); 

    // 4) ?????????? ?????????
    $display("Simulation Finished."); // <-- ???????
    $stop; 
end

endmodule